package simple_uvm_testcase_register_seq_lib_pkg;
    import uvm_pkg::*;
    import autb_csr_agent_pkg::*;
    `include "register_defaults_seq.svh"

    `include "top_on_seq.svh"

endpackage: simple_uvm_testcase_register_seq_lib_pkg