module presistor(.in(a), .out(a));
    inout a;
endmodule
