module presistor(.PLUS(a), .MINUS(a));
    inout a;
endmodule
